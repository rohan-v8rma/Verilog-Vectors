module hello_world; // Name of module same as name of file
    initial
        begin
            $display("Hello World!");
            $finish ;
        end
    endmodule
        